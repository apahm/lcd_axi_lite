`timescale 1 ns / 1 ps

module top_lcd #(
	parameter integer C_S00_AXI_DATA_WIDTH	= 32,
	parameter integer C_S00_AXI_ADDR_WIDTH	= 6
)
(
	input wire  s00_axi_aclk,
	input wire  s00_axi_aresetn,
	input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_awaddr,
	input wire [2 : 0] s00_axi_awprot,
	input wire  s00_axi_awvalid,
	output wire  s00_axi_awready,
	input wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_wdata,
	input wire [(C_S00_AXI_DATA_WIDTH/8)-1 : 0] s00_axi_wstrb,
	input wire  s00_axi_wvalid,
	output wire  s00_axi_wready,
	output wire [1 : 0] s00_axi_bresp,
	output wire  s00_axi_bvalid,
	input wire  s00_axi_bready,
	input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_araddr,
	input wire [2 : 0] s00_axi_arprot,
	input wire  s00_axi_arvalid,
	output wire  s00_axi_arready,
	output wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_rdata,
	output wire [1 : 0] s00_axi_rresp,
	output wire  s00_axi_rvalid,
	input wire  s00_axi_rready,

	// LCD data bus
	output wire [3:0] lcd_data, 
	// LCD: E   (control bit)	
	output wire lcd_e,	
	// LCD: RS  (setup or data)
	output wire lcd_rs,	
	// LCD: R/W (read or write)
	output wire lcd_rw	
);

lcd_control_v1_0_S00_AXI # ( 
	.C_S_AXI_DATA_WIDTH(C_S00_AXI_DATA_WIDTH),
	.C_S_AXI_ADDR_WIDTH(C_S00_AXI_ADDR_WIDTH)
) 
lcd_control_v1_0_S00_AXI_inst 
(
	.S_AXI_ACLK(s00_axi_aclk),
	.S_AXI_ARESETN(s00_axi_aresetn),
	.S_AXI_AWADDR(s00_axi_awaddr),
	.S_AXI_AWPROT(s00_axi_awprot),
	.S_AXI_AWVALID(s00_axi_awvalid),
	.S_AXI_AWREADY(s00_axi_awready),
	.S_AXI_WDATA(s00_axi_wdata),
	.S_AXI_WSTRB(s00_axi_wstrb),
	.S_AXI_WVALID(s00_axi_wvalid),
	.S_AXI_WREADY(s00_axi_wready),
	.S_AXI_BRESP(s00_axi_bresp),
	.S_AXI_BVALID(s00_axi_bvalid),
	.S_AXI_BREADY(s00_axi_bready),
	.S_AXI_ARADDR(s00_axi_araddr),
	.S_AXI_ARPROT(s00_axi_arprot),
	.S_AXI_ARVALID(s00_axi_arvalid),
	.S_AXI_ARREADY(s00_axi_arready),
	.S_AXI_RDATA(s00_axi_rdata),
	.S_AXI_RRESP(s00_axi_rresp),
	.S_AXI_RVALID(s00_axi_rvalid),
	.S_AXI_RREADY(s00_axi_rready),

	.lcd_ready(lcd_ready),
 	.lcd_valid(lcd_valid),
 	.lcd_data_str_0_0(lcd_data_str_0_0),
 	.lcd_data_str_0_1(lcd_data_str_0_1),
 	.lcd_data_str_0_2(lcd_data_str_0_2),
 	.lcd_data_str_0_3(lcd_data_str_0_3),
 	.lcd_data_str_1_0(lcd_data_str_1_0),
 	.lcd_data_str_1_1(lcd_data_str_1_1),
 	.lcd_data_str_1_2(lcd_data_str_1_2),
 	.lcd_data_str_1_3(lcd_data_str_1_3)
);

wire lcd_ready;
wire lcd_valid;
wire [31:0] lcd_data_str_0_0;
wire [31:0] lcd_data_str_0_1;
wire [31:0] lcd_data_str_0_2;
wire [31:0] lcd_data_str_0_3;
wire [31:0] lcd_data_str_1_0;
wire [31:0] lcd_data_str_1_1;
wire [31:0] lcd_data_str_1_2;
wire [31:0] lcd_data_str_1_3;

lcd #(
	.CYCLES_PER_US(50)
)
lcd_inst
(
	.clk(s00_axi_aclk),  
	.rst(~s00_axi_aresetn),  
	.ctrl_lcd({lcd_rs,lcd_rw,lcd_e}),
	.data_lcd(lcd_data),

	.lcd_ready(lcd_ready),
 	.lcd_valid(lcd_valid),
 	.lcd_data_str_0_0(lcd_data_str_0_0),
 	.lcd_data_str_0_1(lcd_data_str_0_1),
 	.lcd_data_str_0_2(lcd_data_str_0_2),
 	.lcd_data_str_0_3(lcd_data_str_0_3),
 	.lcd_data_str_1_0(lcd_data_str_1_0),
 	.lcd_data_str_1_1(lcd_data_str_1_1),
 	.lcd_data_str_1_2(lcd_data_str_1_2),
 	.lcd_data_str_1_3(lcd_data_str_1_3)
);

endmodule
